////////////////////////////////////////////////////////////////////////////////
// Name: Abdelrahman Mohamed
// Course: Digital Verification using SV & UVM (by eng.Kareem Waseem)
//
// Description: FIFO Design (shared package)
// 
////////////////////////////////////////////////////////////////////////////////
package shared_pkg;

//internal signals
    int error_count = 0;
    int correct_count = 0;
    int test_finished = 0;
endpackage